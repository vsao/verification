* SPICE NETLIST
***************************************

.SUBCKT res45 t1 t2
** N=165 EP=2 IP=0 FDC=1
R0 t1 t2 L=2.39774e-05 W=2e-06 $[rnp1] $X=-1525 $Y=-1025 $D=0
.ENDS
***************************************
