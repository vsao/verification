* SPICE NETLIST
***************************************

.SUBCKT resistor_test2 t2 t1
** N=491 EP=2 IP=0 FDC=1
R0 t2 t1 L=0.00018439 W=2e-06 $[rnp1] $X=-1525 $Y=-1025 $D=0
.ENDS
***************************************
