* SPICE NETLIST
***************************************

.SUBCKT pe5_test B S G D
** N=5 EP=4 IP=0 FDC=1
M0 D G S B pe5 L=5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=-235 $Y=-715 $D=0
.ENDS
***************************************
