* SPICE NETLIST
***************************************

.SUBCKT resistor_8strip t1 t2
** N=235 EP=2 IP=0 FDC=1
R0 t1 t2 L=0.00010208 W=2e-06 $[rnp1] $X=-1525 $Y=-1025 $D=0
.ENDS
***************************************
