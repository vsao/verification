* SPICE NETLIST
***************************************

.SUBCKT nwell_res t3 t1 t2
** N=3 EP=3 IP=0 FDC=1
R0 t1 t2 L=1e-05 W=2e-06 $SUB=t3 $[rnw] $X=-1685 $Y=-1145 $D=0
.ENDS
***************************************
