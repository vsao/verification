* SPICE NETLIST
***************************************

.SUBCKT my_resister t2 t1
** N=156 EP=2 IP=0 FDC=1
R0 t2 t1 L=1e-05 W=2e-06 $[rnp1] $X=-1525 $Y=-1025 $D=0
.ENDS
***************************************
