* SPICE NETLIST
***************************************

.SUBCKT ne_test B D G S
** N=4 EP=4 IP=0 FDC=1
M0 S G D B ne L=1.8e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=-1005 $Y=-1395 $D=0
.ENDS
***************************************
