* SPICE NETLIST
***************************************

.SUBCKT cap_test t1 t2
** N=2 EP=2 IP=0 FDC=1
C0 t1 t2 area=4e-10 perimeter=8e-05 $[cmm5t] $X=-1245 $Y=-1245 $D=0
.ENDS
***************************************
